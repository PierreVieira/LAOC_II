library verilog;
use verilog.vl_types.all;
entity p2_mem_ram is
    port(
        clock           : in     vl_logic;
        address         : in     vl_logic_vector(4 downto 0);
        wren            : in     vl_logic;
        data            : in     vl_logic_vector(7 downto 0);
        q               : out    vl_logic_vector(7 downto 0)
    );
end p2_mem_ram;
